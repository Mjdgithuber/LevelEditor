<Level>
<Size width="30" height="30"></Size>
<Tile name="assets\blocks\tree.png" x="0" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="0"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="0"></Tile>
<Tile name="assets\blocks\tree.png" x="9" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="1"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="1"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="1"></Tile>
<Tile name="assets\blocks\tree.png" x="7" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="2"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="2"></Tile>
<Tile name="assets\blocks\tree.png" x="3" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="2"></Tile>
<Tile name="assets\blocks\tree.png" x="6" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="3"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="3"></Tile>
<Tile name="assets\blocks\tree.png" x="3" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="3"></Tile>
<Tile name="assets\blocks\tree.png" x="5" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="4"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="4"></Tile>
<Tile name="assets\blocks\z.png" x="3" y="4"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="5"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="5"></Tile>
<Tile name="assets\blocks\tree.png" x="3" y="5"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="9"></Tile>
<Tile name="assets\blocks\z.png" x="9" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="29"></Tile>
</Level>
