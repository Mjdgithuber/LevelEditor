<Level>
<Size width="150" height="50"></Size>
<Tile name="assets\blocks\grass.png" x="0" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="1"></Tile>
<Tile name="assets\blocks\grass.png" x="1" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="1"></Tile>
<Tile name="assets\blocks\grass.png" x="4" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="1"></Tile>
<Tile name="assets\blocks\grass.png" x="6" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="2"></Tile>
<Tile name="assets\blocks\grass.png" x="1" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="2"></Tile>
<Tile name="assets\blocks\grass.png" x="4" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="3"></Tile>
<Tile name="assets\blocks\grass.png" x="1" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="3"></Tile>
<Tile name="assets\blocks\grass.png" x="7" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="4"></Tile>
<Tile name="assets\blocks\grass.png" x="1" y="4"></Tile>
<Tile name="assets\blocks\grass.png" x="2" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="4"></Tile>
<Tile name="assets\blocks\grass.png" x="4" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="5"></Tile>
<Tile name="assets\blocks\grass.png" x="3" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="5"></Tile>
<Tile name="assets\blocks\grass.png" x="7" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="7"></Tile>
<Tile name="assets\blocks\grass.png" x="2" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="7"></Tile>
<Tile name="assets\blocks\grass.png" x="5" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="7"></Tile>
<Tile name="assets\blocks\grass.png" x="0" y="8"></Tile>
<Tile name="assets\blocks\grass.png" x="1" y="8"></Tile>
<Tile name="assets\blocks\grass.png" x="2" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="8"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="8"></Tile>
<Tile name="assets\blocks\tree.png" x="9" y="8"></Tile>
<Tile name="assets\blocks\tree.png" x="10" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="9"></Tile>
<Tile name="assets\blocks\grass.png" x="5" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="9"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="9"></Tile>
<Tile name="assets\blocks\z.png" x="9" y="9"></Tile>
<Tile name="assets\blocks\tree.png" x="10" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="10"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="10"></Tile>
<Tile name="assets\blocks\tree.png" x="9" y="10"></Tile>
<Tile name="assets\blocks\tree.png" x="10" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="17"></Tile>
<Tile name="assets\blocks\grass.png" x="2" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="19"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="4" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="23"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="2" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="24"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="2" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="25"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="4" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="27"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="2" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="27"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="4" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="28"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="2" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="29"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="7" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="31"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="5" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="32"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="2" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="33"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="2" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="35"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="2" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="36"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="7" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="38"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="2" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="38"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="5" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="39"></Tile>
<Tile name="assets\blocks\treeBorder.png" x="3" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="41"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="41"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="41"></Tile>
<Tile name="assets\blocks\tree.png" x="5" y="41"></Tile>
<Tile name="assets\blocks\tree.png" x="6" y="41"></Tile>
<Tile name="assets\blocks\tree.png" x="7" y="41"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="42"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="42"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="42"></Tile>
<Tile name="assets\blocks\tree.png" x="5" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="43"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="43"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="43"></Tile>
<Tile name="assets\blocks\tree.png" x="5" y="43"></Tile>
<Tile name="assets\blocks\tree.png" x="6" y="43"></Tile>
<Tile name="assets\blocks\tree.png" x="7" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="44"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="44"></Tile>
<Tile name="assets\blocks\z.png" x="3" y="44"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="45"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="45"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="45"></Tile>
<Tile name="assets\blocks\tree.png" x="3" y="45"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="45"></Tile>
<Tile name="assets\blocks\tree.png" x="5" y="45"></Tile>
<Tile name="assets\blocks\tree.png" x="6" y="45"></Tile>
<Tile name="assets\blocks\tree.png" x="7" y="45"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="46"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="46"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="47"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="47"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="48"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="48"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="49"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="49"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="49"></Tile>
<Tile name="assets\blocks\tree.png" x="3" y="49"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="49"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="49"></Tile>
<Building name="assets\buildings\hospital.png" x="5" y="42"></Building>
</Level>
