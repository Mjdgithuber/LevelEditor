<Level>
<Size width="150" height="100"></Size>
<Tile name="assets\blocks\battleSpot_Grass.png" x="0" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="0"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="4" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="0"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="1"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="2"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="1" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="2"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="3"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="4" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="3"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="7" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="3"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="15" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="3"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="29" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="3"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="34" y="3"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="35" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="3"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="4"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="1" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="4"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="24" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="4"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="5"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="2" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="5"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="6"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="5" y="6"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="6" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="6"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="37" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="6"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="7"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="3" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="7"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="32" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="7"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="38" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="7"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="8"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="8"></Tile>
<Tile name="assets\blocks\tree.png" x="9" y="8"></Tile>
<Tile name="assets\blocks\tree.png" x="10" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="8"></Tile>
<Tile name="assets\blocks\battleSpot_Grass.png" x="39" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="8"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="8"></Tile>
<Tile name="assets\blocks\grass.png" x="0" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="9"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="9"></Tile>
<Tile name="assets\blocks\z.png" x="9" y="9"></Tile>
<Tile name="assets\blocks\tree.png" x="10" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="9"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="9"></Tile>
<Tile name="assets\blocks\grass.png" x="0" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="10"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="10"></Tile>
<Tile name="assets\blocks\tree.png" x="9" y="10"></Tile>
<Tile name="assets\blocks\tree.png" x="10" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="10"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="10"></Tile>
<Tile name="assets\blocks\grass.png" x="0" y="11"></Tile>
<Tile name="assets\blocks\grass.png" x="1" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="11"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="12"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="13"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="13"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="14"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="15"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="16"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="17"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="18"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="19"></Tile>
<Tile name="assets\blocks\tree.png" x="3" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="19"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="20"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="21"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="22"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="23"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="23"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="24"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="25"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="26"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="27"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="27"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="28"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="29"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="30"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="31"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="32"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="32"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="33"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="34"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="35"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="36"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="37"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="38"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="38"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="39"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="40"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="41"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="42"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="43"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="44"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="44"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="45"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="46"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="47"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="48"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="49"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="50"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="50"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="51"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="52"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="53"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="54"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="55"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="55"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="56"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="57"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="58"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="59"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="60"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="60"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="61"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="62"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="63"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="64"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="65"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="66"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="66"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="67"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="68"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="69"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="70"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="71"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="72"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="72"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="73"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="74"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="75"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="76"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="76"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="77"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="78"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="79"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="80"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="81"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="81"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="82"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="83"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="84"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="85"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="85"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="86"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="87"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="87"></Tile>
<Tile name="assets\blocks\tree.png" x="0" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="88"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="89"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="90"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="91"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="91"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="92"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="93"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="94"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="95"></Tile>
<Tile name="assets\blocks\tree.png" x="1" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="95"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="96"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="96"></Tile>
<Tile name="assets\blocks\tree.png" x="3" y="96"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="96"></Tile>
<Tile name="assets\blocks\tree.png" x="5" y="96"></Tile>
<Tile name="assets\blocks\tree.png" x="6" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="96"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="96"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="97"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="98"></Tile>
<Tile name="assets\blocks\tree.png" x="2" y="98"></Tile>
<Tile name="assets\blocks\tree.png" x="3" y="98"></Tile>
<Tile name="assets\blocks\tree.png" x="4" y="98"></Tile>
<Tile name="assets\blocks\tree.png" x="5" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="98"></Tile>
<Tile name="assets\blocks\tree.png" x="8" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="74" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="75" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="76" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="77" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="78" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="79" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="80" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="81" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="82" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="83" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="84" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="85" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="86" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="87" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="88" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="89" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="90" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="91" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="92" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="93" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="94" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="95" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="96" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="97" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="98" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="99" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="100" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="101" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="102" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="103" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="104" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="105" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="106" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="107" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="108" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="109" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="110" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="111" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="112" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="113" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="114" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="115" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="116" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="117" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="118" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="119" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="120" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="121" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="122" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="123" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="124" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="125" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="126" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="127" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="128" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="129" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="130" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="131" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="132" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="133" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="134" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="135" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="136" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="137" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="138" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="139" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="140" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="141" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="142" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="143" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="144" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="145" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="146" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="147" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="148" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="149" y="98"></Tile>
<Tile name="assets\blocks\void.png" x="0" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="1" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="2" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="3" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="4" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="5" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="6" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="7" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="8" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="9" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="10" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="11" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="12" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="13" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="14" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="15" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="16" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="17" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="18" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="19" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="20" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="21" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="22" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="23" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="24" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="25" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="26" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="27" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="28" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="29" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="30" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="31" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="32" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="33" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="34" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="35" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="36" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="37" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="38" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="39" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="40" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="41" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="42" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="43" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="44" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="45" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="46" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="47" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="48" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="49" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="50" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="51" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="52" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="53" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="54" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="55" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="56" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="57" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="58" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="59" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="60" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="61" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="62" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="63" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="64" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="65" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="66" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="67" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="68" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="69" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="70" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="71" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="72" y="99"></Tile>
<Tile name="assets\blocks\void.png" x="73" y="99"></Tile>
<Tile name="assets\blocks\void.pn